//////////////////////////////////////////////////////////////////////////////////////////////
 
class mon extends uvm_monitor;
`uvm_component_utils(mon)
 
    uvm_analysis_port#(transaction) send;
    transaction tr;
    virtual spi_i vif;
 
    function new(input string inst = "mon", uvm_component parent = null);
        super.new(inst,parent);
    endfunction
    
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        tr = transaction::type_id::create("tr");
        send = new("send", this);
        if(!uvm_config_db#(virtual spi_i)::get(this,"","vif",vif))//uvm_test_top.env.agent.drv.aif
        `uvm_error("MON","Unable to access Interface");
    endfunction
    
    
    virtual task run_phase(uvm_phase phase);
    forever begin
        @(posedge vif.clk);
        if(vif.rst)
        begin
            tr.op      = rstdut; 
            `uvm_info("MON", "SYSTEM RESET DETECTED", UVM_NONE);
            send.write(tr);
        end
        else if (!vif.rst && vif.wr)
        begin
            @(posedge vif.done);
            tr.op     = writed;
            tr.din    = vif.din;
            tr.addr   = vif.addr;
            tr.err    = vif.err;
            `uvm_info("MON", $sformatf("DATA WRITE addr:%0d data:%0d err:%0d",tr.addr,tr.din,tr.err), UVM_NONE); 
            send.write(tr);
        end
        else if (!vif.rst && !vif.wr)
        begin
            @(posedge vif.done);
            tr.op     = readd; 
            tr.addr   = vif.addr;
            tr.err    = vif.err;
            tr.dout   = vif.dout; 
            `uvm_info("MON", $sformatf("DATA READ addr:%0d data:%0d slverr:%0d",tr.addr,tr.dout,tr.err), UVM_NONE); 
            send.write(tr);
        end
    end
    endtask 
endclass
