// ---------------------------------
//
//
//
//
// ---------------------------------

`ifndef ENV_PKG_SVH
`define ENV_PKG_SVH

 package env_pkg;
 	import uvm_pkg::*;
 	`include "uvm_macros.svh"

	import agent_pkg::*;

	  // Includes:
	`include "sco.svh"
	`include "env.svh"

 endpackage : env_pkg

`endif


