////////////////////////////////////////////////////////////
interface spi_if;
 
    logic clk, rst, cs, miso;
    logic ready, mosi, op_done;
      
endinterface