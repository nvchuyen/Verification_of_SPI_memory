// ----------------------------------
// 31/08/2023
// Nguyen Van Chuyen
//
//
// ----------------------------------


class test_first extends base_test /* base class*/;
	`uvm_component_utils(test_first)

	function new(input string inst, uvm_component c);
		super.new(inst, c);		
	endfunction 


	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		e = 
	endfunction 


endclass : test_first


