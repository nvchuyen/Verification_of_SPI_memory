// ---------------------------------
//
//
//
//
// ---------------------------------

`ifndef SPI_PKG_SVH
`define SPI_PKG_SVH

 package spi_pkg;
 	import uvm_pkg::*;
 	`import "uvm_macros.svh"


 endpackage : spi_pkg

`endif


