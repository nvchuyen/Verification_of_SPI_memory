//
//
// Package Description:
//
package env_pkg;

  // Standard UVM import & include:
import uvm_pkg::*;
`include "uvm_macros.svh"

import agent_pkg::*;


  // Includes:
`include "sco.svh"
`include "env.svh"

endpackage: env_pkg
