//--------------------------------------------
//
//
//
//--------------------------------------------
//
// Class Description
//

package test_lib_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
	
	import env_pkg::*;
	import agent_pkg::*;
	import seq_lib_pkg::*;
	

 // Includes:
`include "test.svh"


endpackage : test_lib_pkg
