
`ifndef SEQ_PKG_SV
`define SEQ_PKG_SV

package seq_lib_pkg;
	
import uvm_pkg::*;
`include "uvm_macros.svh"

	import env_pkg::*;
	import agent_pkg::*;

	`include "transaction.svh"
	`include "read_data.svh"
	`include "read_err.svh"
	`include "reset_dut.svh"
	`include "write_data.svh"
	`include "write_err.svh"
	`include "writeb_readb.svh"


endpackage : seq_lib_pkg
`endif

